module Karatsuba_multipliers_ECC (A,B,C);

    input [7:0] A,B;
    output wire [15:0] C;

    wire [7:0] M [0:7];

    assign M[0][0] = A[0] & B[0];
    assign M[1][0] = A[1] & B[1];
    assign M[2][0] = A[2] & B[2];
    assign M[3][0] = A[3] & B[3];
    assign M[4][0] = A[4] & B[4];
    assign M[5][0] = A[5] & B[5];
    assign M[6][0] = A[6] & B[6];
    assign M[7][0] = A[7] & B[7];
    assign M[0][1] = (A[0] ^ A[1]) & (B[0] ^ B[1]);
    assign M[0][2] = (A[0] ^ A[2]) & (B[0] ^ B[2]);
    assign M[0][3] = (A[0] ^ A[3]) & (B[0] ^ B[3]);
    assign M[0][4] = (A[0] ^ A[4]) & (B[0] ^ B[4]);
    assign M[0][5] = (A[0] ^ A[5]) & (B[0] ^ B[5]);
    assign M[0][6] = (A[0] ^ A[6]) & (B[0] ^ B[6]);
    assign M[0][7] = (A[0] ^ A[7]) & (B[0] ^ B[7]);
    assign M[1][2] = (A[1] ^ A[2]) & (B[1] ^ B[2]);
    assign M[1][3] = (A[1] ^ A[3]) & (B[1] ^ B[3]);
    assign M[1][4] = (A[1] ^ A[4]) & (B[1] ^ B[4]);
    assign M[1][5] = (A[1] ^ A[5]) & (B[1] ^ B[5]);
    assign M[1][6] = (A[1] ^ A[6]) & (B[1] ^ B[6]);
    assign M[1][7] = (A[1] ^ A[7]) & (B[1] ^ B[7]);
    assign M[2][3] = (A[2] ^ A[3]) & (B[2] ^ B[3]);
    assign M[2][4] = (A[2] ^ A[4]) & (B[2] ^ B[4]);
    assign M[2][5] = (A[2] ^ A[5]) & (B[2] ^ B[5]);
    assign M[2][6] = (A[2] ^ A[6]) & (B[2] ^ B[6]);
    assign M[2][7] = (A[2] ^ A[7]) & (B[2] ^ B[7]);
    assign M[3][4] = (A[3] ^ A[4]) & (B[3] ^ B[4]);
    assign M[3][5] = (A[3] ^ A[5]) & (B[3] ^ B[5]);
    assign M[3][6] = (A[3] ^ A[6]) & (B[3] ^ B[6]);
    assign M[3][7] = (A[3] ^ A[7]) & (B[3] ^ B[7]);
    assign M[4][5] = (A[4] ^ A[5]) & (B[4] ^ B[5]);
    assign M[4][6] = (A[4] ^ A[6]) & (B[4] ^ B[6]);
    assign M[4][7] = (A[4] ^ A[7]) & (B[4] ^ B[7]);
    assign M[5][6] = (A[5] ^ A[6]) & (B[5] ^ B[6]);
    assign M[5][7] = (A[5] ^ A[7]) & (B[5] ^ B[7]);
    assign M[6][7] = (A[6] ^ A[7]) & (B[6] ^ B[7]);
    assign C[0] = M[0][0];
    assign C[1] = M[0][1] ^ M[0][0] ^ M[1][0];
    assign C[2] = M[0][2] ^ M[0][0] ^ M[1][0] ^ M[2][0];
    assign C[3] = M[0][3] ^ M[1][2] ^ M[0][0] ^ M[1][0] ^ M[2][0] ^ M[3][0];
    assign C[4] = M[0][4] ^ M[1][3] ^ M[0][0] ^ M[1][0] ^ M[2][0] ^ M[3][0] ^ M[4][0];
    assign C[5] = M[0][5] ^ M[1][4] ^ M[2][3] ^ M[0][0] ^ M[1][0] ^ M[2][0] ^ M[3][0] ^ M[4][0] ^ M[5][0];
    assign C[6] = M[0][6] ^ M[1][5] ^ M[2][4] ^ M[0][0] ^ M[1][0] ^ M[2][0] ^ M[3][0] ^ M[4][0] ^ M[5][0] ^ M[6][0];
    assign C[7] = M[0][7] ^ M[1][6] ^ M[2][5] ^ M[3][4] ^ M[0][0] ^ M[1][0] ^ M[2][0] ^ M[3][0] ^ M[4][0] ^ M[5][0] ^ M[6][0] ^ M[7][0];
    assign C[8] = M[1][7] ^ M[2][6] ^ M[3][5] ^ M[1][0] ^ M[2][0] ^ M[3][0] ^ M[4][0] ^ M[5][0] ^ M[6][0] ^ M[7][0];
    assign C[9] = M[2][7] ^ M[3][6] ^ M[4][5] ^ M[2][0] ^ M[3][0] ^ M[4][0] ^ M[5][0] ^ M[6][0] ^ M[7][0];
    assign C[10] = M[3][7] ^ M[4][6] ^ M[3][0] ^ M[4][0] ^ M[5][0] ^ M[6][0] ^ M[7][0];
    assign C[11] = M[4][7] ^ M[5][6] ^ M[4][0] ^ M[5][0] ^ M[6][0] ^ M[7][0];
    assign C[12] = M[5][7] ^ M[5][0] ^ M[6][0] ^ M[7][0];
    assign C[13] = M[6][7] ^ M[6][0] ^ M[7][0];
    assign C[14] = M[7][0];
    assign C[15] = 0;   
    
endmodule